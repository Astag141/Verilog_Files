module mealy_seq_detector (
    input clk,
    input reset,
    input x,
    output reg z
);
    typedef enum logic [1:0] {
        S0, S1, S2, S3
    } state_t;

    state_t current_state, next_state;

    always @(posedge clk or posedge reset) begin
        if (reset)
            current_state <= S0;
        else
            current_state <= next_state;
    end

    always @(*) begin
        z = 0;
        case (current_state)
            S0: next_state = (x == 1) ? S1 : S0;
            S1: next_state = (x == 0) ? S2 : S1;
            S2: next_state = (x == 1) ? S3 : S0;
            S3: begin
                if (x == 1) begin
                    next_state = S1;
                    z = 1;
                end else begin
                    next_state = S2;
                    z = 0;
                end
            end
        endcase
    end
endmodule