module tb_parity_generator; reg [3:0] data; wire parity; parity_generator uut (.data(data), .parity(parity)); initial begin data=4'b1010; #5 $display("Data=%b Parity=%b", data, parity); end endmodule