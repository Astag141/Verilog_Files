module tb_half_subtractor;
    reg a, b;
    wire diff, borrow;
    half_subtractor uut (.a(a), .b(b), .diff(diff), .borrow(borrow));
    initial begin
        a=0; b=0; #10;
        a=0; b=1; #10;
        a=1; b=0; #10;
        a=1; b=1; #10;
        $finish;
    end
initial $monitor("tb_a=%b tb_b=%b tb_diff=%b tb_borrow=%b",a,b,diff,borrow);
endmodule
