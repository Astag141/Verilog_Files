module lut4x1(input [3:0] addr, output y); assign y = (addr == 4'b0000) ? 1'b0 : (addr == 4'b0001) ? 1'b1 : (addr == 4'b0010) ? 1'b0 : (addr == 4'b0011) ? 1'b1 : (addr == 4'b0100) ? 1'b1 : (addr == 4'b0101) ? 1'b0 : (addr == 4'b0110) ? 1'b1 : (addr == 4'b0111) ? 1'b0 : (addr == 4'b1000) ? 1'b0 : (addr == 4'b1001) ? 1'b1 : 1'b0; endmodule