module encoder2x1(input [1:0] in, output y);
  assign y = in[1];
endmodule

